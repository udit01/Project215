--Created By:-
--Shashwat Shivam & Udit Jain
--2016CS10328 & 2016CS10327



----------------------------------------------------------------------------------
-- Company:
-- Engineer:
--
-- Create Date: 27.08.2017 08:20:05
-- Design Name:
-- Module Name: display - struc
-- Project Name:
-- Target Devices:
-- Tool Versions:
-- Description:
--
-- Dependencies:
--
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity uart_tx is
PORT (
  data_input:in std_logic_vector(15 downto 0):="0000000000000000";
  clk:in std_logic;
  reset:in STD_LOGIC:='0';--upButton
  send:in STD_LOGIC:='0';--middle button
  sendL:in std_logic:='0';
  sendR:in std_logic:='0';
  data:out STD_LOGIC;--RS32
  sim_mode:in std_logic;--down Button
--  busy:out std_logic;
  led:out std_logic_vector(15 downto 0);
  cathode:out std_logic_vector(6 downto 0);
  anode:out std_logic_vector(3 downto 0)
  --to leds?
	);

end uart_tx;

architecture structural of uart_tx is
  -- COMPONENT display is
  --   port(
  --   data: in std_logic_vector(15 downto 0);
  -- 	clk: in std_logic;
  --   sim_mode: in std_logic;
  -- 	anode : out std_logic_vector (3 downto 0);
  -- 	cathode : OUT std_logic_vector (6 downto 0)
  --   )
  -- END COMPONENT;

signal sending_pos : integer :=0;
signal loop_number : integer :=69;
signal loop_number2 : integer :=897;
signal data_internal,final_clock,comparator1,comparator2,general_comparator,general_comparator2: std_logic:='1';
signal busy_internal,busy_internal1,busy_internal2,busy_internal3,send_pulse,send_pulseL,send_pulseR,clock: std_logic:='0';
signal counter: std_logic_vector(8 downto 0):="000000000";
signal data1,data2:std_logic_vector(7 downto 0):="00000000";

type t_Memory is array (0 to 69) of std_logic_vector(7 downto 0);
signal data_arr : t_Memory:=
("00001101","00001010","01010000","01110010","01101111","01101010","01100101","01100011","01110100","00100000","01000010","01111001","00111010","00101101","00001101","00001010","01010011","01101000","01100001","01110011","01101000","01110111","01100001","01110100","00100000","01010011","01101000","01101001","01110110","01100001","01101101","00001101","00001010","00110010","00110000","00110001","00110110","01000011","01010011","00110001","00110000","00110011","00110010","00111000","00001101","00001010","01010101","01100100","01101001","01110100","00100000","01001010","01100001","01101001","01101110","00001101","00001010","00110010","00110000","00110001","00110110","01000011","01010011","00110001","00110000","00110011","00110010","00110111","00001101","00001010");

type t_Memory2 is array (0 to 897) of std_logic_vector(7 downto 0);
signal data_arr2 : t_Memory2:=("00001101","00001010","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00101000","00100000","00100000","00101001","00100000","00101000","01000000","01000000","00101001","00100000","00101000","00100000","00101001","00100000","00100000","00101000","01000000","00101001","00100000","00100000","00101000","00101001","00100000","00100000","00100000","00100000","01000000","01000000","00100000","00100000","00100000","00100000","01001111","00100000","00100000","00100000","00100000","00100000","01000000","00100000","00100000","00100000","00100000","00100000","01001111","00100000","00100000","00100000","00100000","00100000","01000000","00001101","00001010","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00101000","01000000","01000000","01000000","00101001","00001101","00001010","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00101000","00100000","00100000","00100000","00100000","00101001","00001101","00001010","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00101000","01000000","01000000","01000000","01000000","00101001","00001101","00001010","00001101","00001010","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00101000","00100000","00100000","00100000","00101001","00001101","00001010","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00111101","00111101","00111101","00111101","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","00001101","00001010","00100000","00100000","00100000","00100000","01011111","01000100","00100000","01011111","01111100","00100000","00100000","01111100","01011111","01011111","01011111","01011111","01011111","01011111","01011111","00101111","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","01011100","01011111","01011111","01001001","01011111","01001001","01011111","01011111","01011111","01011111","01011111","00111101","00111101","00111101","01011111","01011111","01111100","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01111100","00001101","00001010","00100000","00100000","00100000","00100000","00100000","01111100","00101000","01011111","00101001","00101101","00101101","00101101","00100000","00100000","01111100","00100000","00100000","00100000","01001000","01011100","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","00101111","00100000","01111100","00100000","00100000","00100000","01111100","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00111101","01111100","01011111","01011111","01011111","00100000","01011111","01011111","01011111","01111100","00100000","00100000","00100000","00100000","00100000","00100000","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","00001101","00001010","00100000","00100000","00100000","00100000","00100000","00101111","00100000","00100000","00100000","00100000","00100000","01111100","00100000","00100000","01111100","00100000","00100000","00100000","01001000","00100000","00100000","01111100","00100000","00100000","01111100","00100000","00100000","00100000","00100000","00100000","01111100","00100000","00100000","00100000","01111100","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","01111100","01111100","01011111","01111100","00100000","01111100","01011111","01111100","01111100","00100000","00100000","00100000","00100000","00100000","01011111","01111100","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","01011100","01011111","01011111","01011111","00001101","00001010","00100000","00100000","00100000","00100000","01111100","00100000","00100000","00100000","00100000","00100000","00100000","01111100","00100000","00100000","01111100","00100000","00100000","00100000","01001000","00100000","00100000","01111100","01011111","01011111","00101101","00101101","00101101","00101101","00101101","00101101","00101101","00101101","00101101","00101101","00101101","00101101","00101101","00101101","00101101","00101101","00101101","00101101","00101101","00101101","01111100","00100000","01011011","01011111","01011111","01011111","01011101","00100000","01111100","00100000","00100000","00100000","00111101","01111100","00001101","00001010","00100000","00100000","00100000","00100000","01111100","00100000","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01111100","01011111","01011111","01011111","01001000","01011111","01011111","00101111","01011111","01011111","01111100","01011111","01011111","01011111","01011111","01011111","00101111","01011011","01011101","01011011","01011101","01111110","01011100","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01111100","00100000","00100000","00100000","00100000","00100000","00100000","00100000","01111100","00100000","00100000","00100000","00101101","01111100","00001101","00001010","00100000","00100000","00100000","00100000","01111100","00101111","00100000","01111100","00100000","00100000","00100000","01111100","00101101","00101101","00101101","00101101","00101101","00101101","00101101","00101101","00101101","00101101","00101101","01001001","01011111","01011111","01011111","01011111","01011111","01001001","00100000","01011011","01011101","01011011","01011101","00100000","01011011","01011101","00100000","00100000","01000100","00100000","00100000","00100000","01111100","00111101","00111101","00111101","00111101","00111101","00111101","00111101","01111100","01011111","01011111","01011111","01011111","01111100","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","00001101","00001010","00100000","00100000","01011111","01011111","00101111","00100000","00111101","01111100","00100000","01101111","00100000","01111100","00111101","00101101","01111110","01111110","01011100","00100000","00100000","00101111","01111110","01111110","01011100","00100000","00100000","00101111","01111110","01111110","01011100","00100000","00100000","00101111","01111110","01111110","01011100","00100000","01011111","01011111","01011111","01011111","01011001","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01111100","01011111","01011111","01111100","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","01011111","00001101","00001010","00100000","00100000","00100000","01111100","00101111","00101101","00111101","01111100","01011111","01011111","01011111","01111100","00111101","01001111","00111101","00111101","00111101","00111101","00111101","01001111","00111101","00111101","00111101","00111101","00111101","01001111","00111101","00111101","00111101","00111101","00111101","01001111","00100000","00100000","00100000","01111100","01011111","01011111","01011111","01011111","01011111","00101111","01111110","01011100","01011111","01011111","01011111","00101111","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","01111100","01011111","01000100","01011111","01011111","01000100","01011111","01011111","01000100","01011111","01111100","00100000","00100000","01111100","01011111","01000100","01011111","01011111","01000100","01011111","01011111","01000100","00001101","00001010","00100000","00100000","00100000","00100000","01011100","01011111","00101111","00100000","00100000","00100000","00100000","00100000","00100000","01011100","01011111","01011111","00101111","00100000","00100000","01011100","01011111","01011111","00101111","00100000","00100000","01011100","01011111","01011111","00101111","00100000","00100000","01011100","01011111","01011111","00101111","00100000","00100000","00100000","00100000","00100000","00100000","01011100","01011111","00101111","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","00100000","01011100","01011111","00101111","00100000","00100000","00100000","01011100","01011111","00101111","00100000","00100000","00100000","00100000","01011100","01011111","00101111","00100000","00100000","00100000","01011100","00001101","00001010");

begin



data1<=data_input(15 downto 8);
data2<=data_input(7 downto 0);

comparator1<= '1' when not((data1 and counter(7 downto 0)) =  "00000000" )
--comparator1<= '1' when not(("01000000" and counter(7 downto 0)) =  "00000000" )
                else '0';

comparator2<= '1' when not((data2 and counter(7 downto 0)) =  "00000000" )
--comparator2<= '1' when not(("01000000" and counter(7 downto 0)) =  "00000000" )
                else '0';

general_comparator<='1' when not((data_arr(sending_pos) and counter(7 downto 0)) =  "00000000" )
--comparator2<= '1' when not(("01000000" and counter(7 downto 0)) =  "00000000" )
                else '0';

 general_comparator2<='1' when not((data_arr2(sending_pos) and counter(7 downto 0)) =  "00000000" )
                --comparator2<= '1' when not(("01000000" and counter(7 downto 0)) =  "00000000" )
                                else '0';

--led(14 downto 1)<= data_input(14 downto 1);
--led(0)<= data_internal;
--led(15)<= data_internal;
led <= data_input;

final_clock<= clk when sim_mode='1' else clock;

ssd:ENTITY WORK.display(struc)
  PORT MAP(data_input=>data_input,clk=>clk,sim_mode=>sim_mode,anode=>anode,cathode=>cathode);

clocker: ENTITY WORK.transmitter_clock(struc)
	PORT MAP(clock=>clk,out_clock=>clock);


pulse: ENTITY WORK.level2pulseConverter(struc)
PORT MAP(clk=>final_clock,in1=>send,out1=>send_pulse);

pulse2: ENTITY WORK.level2pulseConverter(struc)
PORT MAP(clk=>final_clock,in1=>sendL,out1=>send_pulseL);
pulse3: ENTITY WORK.level2pulseConverter(struc)
PORT MAP(clk=>final_clock,in1=>sendR,out1=>send_pulseR);

--    send_pulse <= send;
--	display: ENTITY WORK.display(struc)
--	PORT MAP(clk=>clk,data=>data_input,anode=>anode,cathode=>cathode);

data<=data_internal;
--busy<=busy_internal;
busy_internal<=busy_internal1 or busy_internal2 or busy_internal3;
process(final_clock,reset)
begin
    if(reset='1') then

                        data_internal<='1';
                        busy_internal1<='0';
                        busy_internal2<='0';
                        busy_internal3<='0';
                        counter<="000000000";
                        sending_pos<=0;

    elsif (rising_edge(final_clock)) then

                        if(send_pulse='1' and busy_internal='0') then

                                                   busy_internal1<='1';
                                                   data_internal<='0';
                                                   counter<="000000001";
                                                   sending_pos<=0;

                        elsif(send_pulseL='1' and busy_internal='0') then

                                                    busy_internal2<='1';
                                                    data_internal<='0';
                                                   counter<="000000001";
                                                   sending_pos<=0;

                           elsif(send_pulseR='1' and busy_internal='0') then

                                                   busy_internal3<='1';
                                                   data_internal<='0';
                                                  counter<="000000001";
                                                  sending_pos<=0;

                        elsif(busy_internal1='1') then
                                                  if(counter="100000000") then

                                                                    data_internal<='1';
                                                                    counter<="000000000";

                                                                    if(sending_pos=0) then
                                                                        sending_pos<=1;
--                                                                        counter<="000000000";
                                                                    else
                                                                    busy_internal1<='0';
                                                                    sending_pos<=0;
                                                                    end if;

                                                    elsif(sending_pos=0)       then
--                                                                   elsif((data1 or counter(7 downto 0))> "00000000") then
                                                                        data_internal<=comparator1;
--                                                                    else
--                                                                        data_internal<='0';
--                                                                    end if;
                                                                    counter<=counter(7 downto 0) & '0';
                                                     else
--                                                                    if((data2 or counter(7 downto 0))> "00000000") then
                                                                     if(counter="000000000") then
                                                                                        data_internal<='0';
                                                                                     counter<="000000001";
--                                                                        sending_pos<='0';
                                                                      else
                                                                                    data_internal<=comparator2;
                                                                                    counter<=counter(7 downto 0) & '0';
                                                                      end if;
--                                                                    else
--                                                                        data_internal<='0';
--                                                                    end if;
                                                      end if;
                               elsif(busy_internal2='1') then
                                                               if(counter="100000000") then
                                                                                 data_internal<='1';
                                                                                 counter<="000000000";
                                                                                 if(sending_pos=loop_number) then
                                                                                    busy_internal2<='0';
                                                                                     sending_pos<=0;
                                                                                 else
                                                                                  sending_pos<=sending_pos+1;
                                                                                 end if;
                                                                  else
                                                                                  if(counter="000000000") then
                                                                                                     data_internal<='0';
                                                                                                  counter<="000000001";
                                                                                   else
                                                                                                 data_internal<=general_comparator;
                                                                                                 counter<=counter(7 downto 0) & '0';
                                                                                   end if;
                                                                   end if;
                             elsif(busy_internal3='1') then
                                                             if(counter="100000000") then
                                                                               data_internal<='1';
                                                                               counter<="000000000";
                                                                               if(sending_pos=loop_number2) then
                                                                                  busy_internal3<='0';
                                                                                   sending_pos<=0;
                                                                               else
                                                                                sending_pos<=sending_pos+1;
                                                                               end if;
                                                                else
                                                                                if(counter="000000000") then
                                                                                                   data_internal<='0';
                                                                                                counter<="000000001";
                                                                                 else
                                                                                               data_internal<=general_comparator2;
                                                                                               counter<=counter(7 downto 0) & '0';
                                                                                 end if;
                                                                 end if;

                            end if;

            end if;
--    end if;
end process;



end structural;
